* Ring Oscillator test circuit for Standard Cell Characterization
.option scale=1E-6

* Include the SkyWater Standard Cells
.include /data02/ECE4203/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

* Include SkyWater sky130 device models
.lib "/data02/ECE4203/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

.temp TEMPVALUE
.param cpar=CPARVALUE
.param fanout=FANOUTVALUE

* Subcircuit "testcell" contains the standard cell we are testing.
* 
*  Replace "sky130_fd_sc_hd__nand2_2" with a different cell as desired.
*
*  Note that the other inputs to the gate being tested should be connected to 
*   pull_up or pull_down, in order the make sure the gate will switch.
*
.subckt testcell in out pwr gnd
R1 pull_up pwr 0 
R2 pull_down gnd 0 
X1 CELLINPUTSVALUE gnd gnd pwr pwr out sky130_fd_sc_hd__CELLNAMEVALUE
.ends 

* Subcircuit "fanoutload" creates additional fanout loading, from +0 to +5
*  note that the fanout is already 1 in the ring oscillator
* 
.subckt fanoutload in pwr gnd
.if (fanout==1)
Cempty in 0 0.001f
.elseif (fanout==2)
X1 in uc1 pwr gnd testcell
.elseif (fanout==3)
X1 in uc1 pwr gnd testcell
X2 in uc2 pwr gnd testcell
.elseif (fanout==4)
X1 in uc1 pwr gnd testcell
X2 in uc2 pwr gnd testcell
X3 in uc3 pwr gnd testcell
.elseif (fanout==5)
X1 in uc1 pwr gnd testcell
X2 in uc2 pwr gnd testcell
X3 in uc3 pwr gnd testcell
X4 in uc4 pwr gnd testcell
.elseif (fanout==6)
X1 in uc1 pwr gnd testcell
X2 in uc2 pwr gnd testcell
X3 in uc3 pwr gnd testcell
X4 in uc4 pwr gnd testcell
X5 in uc5 pwr gnd testcell
.endif
.ends

X1 out11 out1 VPWR VGND testcell
C1 out1 0 C='cpar'
X1fan out1 VPWR VGND fanoutload

X2 out1 out2 VPWR VGND testcell
C2 out2 0 C='cpar'
X2fan out2 VPWR VGND fanoutload

X3 out2 out3 VPWR VGND testcell
C3 out3 0 C='cpar'
X3fan out3 VPWR VGND fanoutload

X4 out3 out4 VPWR VGND testcell
C4 out4 0 C='cpar'
X4fan out4 VPWR VGND fanoutload

X5 out4 out5 VPWR VGND testcell
C5 out5 0 C='cpar'
X5fan out5 VPWR VGND fanoutload

X6 out5 out6 VPWR VGND testcell
C6 out6 0 C='cpar'
X6fan out6 VPWR VGND fanoutload

X7 out6 out7 VPWR VGND testcell
C7 out7 0 C='cpar'
X7fan out7 VPWR VGND fanoutload

X8 out7 out8 VPWR VGND testcell
C8 out8 0 C='cpar'
X8fan out8 VPWR VGND fanoutload

X9 out8 out9 VPWR VGND testcell
C9 out9 0 C='cpar'
X9fan out9 VPWR VGND fanoutload

X10 out9 out10 VPWR VGND testcell
C10 out10 0 C='cpar'
X10fan out10 VPWR VGND fanoutload

X11 out10 out11 VPWR VGND testcell
C11 out11 0 C='cpar'
X11fan out11 VPWR VGND fanoutload

I1 out1 0 PULSE 0 0.1u 1e-9 0.1e-9 0.1e-9 1e-9 100e-6

VDD VPWR 0 1.8
VSS VGND 0 0

.control
    tran 10p 30n 
    meas tran period TRIG v(out11) td=15n VAL=0.9 RISE=1 TARG v(out11) td=15n VAL=0.9 RISE=2
    meas tran tpd_rise TRIG v(out10) td=15n VAL=0.9 FALL=1 TARG v(out11) td=15n VAL=0.9 RISE=1
    meas tran tpd_fall TRIG v(out10) td=15n VAL=0.9 RISE=1 TARG v(out11) td=15n VAL=0.9 FALL=1
    plot v(out10) v(out11) 
.endc

.end
